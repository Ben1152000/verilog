module alu (
    input wire [2:0] op
,   input wire [31:0] in1
,   input wire [31:0] in2
,   output reg [31:0] out  /* don't forget to add flags */
);

    always @* begin
        case (op)
            3'b000: out = in1 & in2;  /* and */
            3'b001: out = in1 | in2;  /* or  */
            3'b010: out = in1 + in2;  /* add */
            3'b011: out = 32'h0;
            3'b100: out = 32'h0;
            3'b101: out = 32'h0;
            3'b110: out = in1 - in2;  /* sub */
            3'b111: out = in1 < in2;  /* slt */
        endcase
    end

endmodule
